`timescale 1ns / 1ps

module RF(
    );


endmodule
